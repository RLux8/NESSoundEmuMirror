--
-- VHDL Architecture audiotest_lib.pulseTBctrl.behav
--
-- Created:
--          by - redacted.redacted (pc025)
--          at - 15:44:50 01/08/24
--
-- using Mentor Graphics HDL Designer(TM) 2022.3 Built on 14 Jul 2022 at 13:56:12
--
LIBRARY ieee;
USE IEEE.numeric_std.all;
use ieee.std_logic_1164.all;

ARCHITECTURE behav OF pulseTBctrl IS
  type stateT is (INIT, WRITE1, WRITE2, WRITE3, WRITE4, WRITE5, DONE);
  signal state: stateT;
BEGIN
  fsm_transitions : process(clk, res_n) is
    variable state_int: stateT;
  begin
    if res_n = '0' then
      state_int := INIT;
    else
      if clk'event and clk = '1' then
        if apuclk then
          case state_int is
          when INIT => state_int := WRITE1;
          when WRITE1 => state_int := WRITE2;
          when WRITE2 => state_int := WRITE3;
          when WRITE3 => state_int := WRITE4;
          when WRITE4 => state_int := WRITE5; 
          when WRITE5 => state_int := DONE;
          when DONE => null;
          end case;
        end if;
      end if;
    end if;
    
    state <= state_int;
  end process fsm_transitions;
  
  fsm_outputs: process(state) is
  begin
    case state is
      when INIT => 
        addr <= (false, false);
        data <=  (others => false);
        wr <= false;
      when WRITE1 =>
        addr <= (false, false);
        data <=  (false, false, true, true, true, true, true, true);
        wr <= true;
      when WRITE2 =>
        addr <= (false,true);
        data <= (true, false, false, true, false, false, false, true);
        wr <= true;
      
      when WRITE3 =>
        addr <= (true, false);
        data <= (others => true);
        wr <= true;
    
      when WRITE4 =>
        addr <= (true, true);
        data <= (3 => true, others => false); --B"01011000";
        wr <= true;
       
      when WRITE5 =>
        addr <= (false, false);
        data <=  (false, false, false, false, false, false, true, true);
        wr <= true; 
      
      when DONE => wr <= false;
    end case;
    mode <= false;
    genint <= false;
    resctr <= false;
  end process fsm_outputs;
END ARCHITECTURE behav;