--
-- VHDL Entity audiotest_lib.clk_res_gen.arch_name
--
-- Created:
--          by - redacted.redacted (pc038)
--          at - 14:28:32 12/13/23
--
-- using Mentor Graphics HDL Designer(TM) 2022.3 Built on 14 Jul 2022 at 13:56:12
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
entity clk_res_gen is
port(
clk: out std_logic;
res_n: out std_logic
);
end entity clk_res_gen;


